library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;


entity Top_tb is
end Top_tb;


architecture top_basys_tb of Top_tb is
begin



end top_basys_tb;

